library verilog;
use verilog.vl_types.all;
entity COTROL_CIRCUIT_vlg_vec_tst is
end COTROL_CIRCUIT_vlg_vec_tst;
