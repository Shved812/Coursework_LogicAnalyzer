library verilog;
use verilog.vl_types.all;
entity EDGE_CODER_vlg_vec_tst is
end EDGE_CODER_vlg_vec_tst;
