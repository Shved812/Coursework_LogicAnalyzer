library verilog;
use verilog.vl_types.all;
entity modulator_vlg_check_tst is
    port(
        \out\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end modulator_vlg_check_tst;
