library verilog;
use verilog.vl_types.all;
entity valider_vlg_vec_tst is
end valider_vlg_vec_tst;
