library verilog;
use verilog.vl_types.all;
entity modulator_vlg_vec_tst is
end modulator_vlg_vec_tst;
