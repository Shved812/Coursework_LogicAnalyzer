library verilog;
use verilog.vl_types.all;
entity ARCHIVATOR_vlg_vec_tst is
end ARCHIVATOR_vlg_vec_tst;
