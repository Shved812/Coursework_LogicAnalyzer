library verilog;
use verilog.vl_types.all;
entity sender_counter_vlg_vec_tst is
end sender_counter_vlg_vec_tst;
