library verilog;
use verilog.vl_types.all;
entity counter_locked_vlg_check_tst is
    port(
        clk_out         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end counter_locked_vlg_check_tst;
