library verilog;
use verilog.vl_types.all;
entity parallelizer_vlg_vec_tst is
end parallelizer_vlg_vec_tst;
