library verilog;
use verilog.vl_types.all;
entity counter_locked_vlg_vec_tst is
end counter_locked_vlg_vec_tst;
