library verilog;
use verilog.vl_types.all;
entity valider_vlg_check_tst is
    port(
        switch          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end valider_vlg_check_tst;
